


module top #(
    parameter ADDR_WIDTH = 32,
    parameter DATA_WIDTH = 32
) (
    input  logic clk_i,
    input  logic rst_ni

    // Instructions
    // input  logic instr_data_i
);

    import toothless_pkg::*;


endmodule
